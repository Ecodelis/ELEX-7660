// File: upDownCount.sv
// Description: Simple state machine that counts up or down 
//              based on the input signal upDown.
// Author: Marcus Fu
// Date: 2025-01-17

module upDownCnt3 ( input logic upDown
                    output logic [2:0] count,
                    input logic clk) ;


endmodule